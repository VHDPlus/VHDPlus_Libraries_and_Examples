-- LogicAnalyzer.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LogicAnalyzer is
	port (
		acq_clk        : in std_logic                     := '0';             -- acq_clk.clk
		acq_data_in    : in std_logic_vector(31 downto 0) := (others => '0'); --     tap.acq_data_in
		acq_trigger_in : in std_logic_vector(0 downto 0)  := (others => '0')  --        .acq_trigger_in
	);
end entity LogicAnalyzer;

architecture rtl of LogicAnalyzer is
	component sld_signaltap is
		generic (
			sld_data_bits               : integer := 1;
			sld_sample_depth            : integer := 128;
			sld_ram_block_type          : string  := "AUTO";
			sld_storage_qualifier_mode  : string  := "OFF";
			sld_trigger_bits            : integer := 1;
			sld_trigger_level           : integer := 1;
			sld_trigger_in_enabled      : integer := 0;
			sld_enable_advanced_trigger : integer := 0;
			sld_trigger_level_pipeline  : integer := 1;
			sld_trigger_pipeline        : integer := 0;
			sld_ram_pipeline            : integer := 0;
			sld_counter_pipeline        : integer := 0;
			sld_node_info               : integer := 806383104;
			sld_incremental_routing     : integer := 0;
			sld_node_crc_bits           : integer := 32;
			sld_node_crc_hiword         : integer := 12345;
			sld_node_crc_loword         : integer := 19899
		);
		port (
			acq_data_in    : in std_logic_vector(31 downto 0) := (others => 'X'); -- acq_data_in
			acq_trigger_in : in std_logic_vector(0 downto 0)  := (others => 'X'); -- acq_trigger_in
			acq_clk        : in std_logic                     := 'X'              -- clk
		);
	end component sld_signaltap;

begin

	signaltap_ii_logic_analyzer_0 : component sld_signaltap
		generic map (
			sld_data_bits               => 32,
			sld_sample_depth            => 256,
			sld_ram_block_type          => "AUTO",
			sld_storage_qualifier_mode  => "OFF",
			sld_trigger_bits            => 1,
			sld_trigger_level           => 1,
			sld_trigger_in_enabled      => 0,
			sld_enable_advanced_trigger => 0,
			sld_trigger_level_pipeline  => 1,
			sld_trigger_pipeline        => 0,
			sld_ram_pipeline            => 0,
			sld_counter_pipeline        => 0,
			sld_node_info               => 806383104,
			sld_incremental_routing     => 0,
			sld_node_crc_bits           => 32,
			sld_node_crc_hiword         => 19939,
			sld_node_crc_loword         => 16463
		)
		port map (
			acq_data_in    => acq_data_in,    --     tap.acq_data_in
			acq_trigger_in => acq_trigger_in, --        .acq_trigger_in
			acq_clk        => acq_clk         -- acq_clk.clk
		);

end architecture rtl; -- of LogicAnalyzer
