-- megafunction wizard: %Triple-Speed Ethernet Intel FPGA IP v18.1%
-- GENERATION: XML
-- Ethernet.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Ethernet is
	port (
		clk           : in  std_logic                     := '0';             -- control_port_clock_connection.clk
		reset         : in  std_logic                     := '0';             --              reset_connection.reset
		reg_addr      : in  std_logic_vector(7 downto 0)  := (others => '0'); --                  control_port.address
		reg_data_out  : out std_logic_vector(31 downto 0);                    --                              .readdata
		reg_rd        : in  std_logic                     := '0';             --                              .read
		reg_data_in   : in  std_logic_vector(31 downto 0) := (others => '0'); --                              .writedata
		reg_wr        : in  std_logic                     := '0';             --                              .write
		reg_busy      : out std_logic;                                        --                              .waitrequest
		tx_clk        : in  std_logic                     := '0';             --   pcs_mac_tx_clock_connection.clk
		rx_clk        : in  std_logic                     := '0';             --   pcs_mac_rx_clock_connection.clk
		set_10        : in  std_logic                     := '0';             --         mac_status_connection.set_10
		set_1000      : in  std_logic                     := '0';             --                              .set_1000
		eth_mode      : out std_logic;                                        --                              .eth_mode
		ena_10        : out std_logic;                                        --                              .ena_10
		m_rx_d        : in  std_logic_vector(3 downto 0)  := (others => '0'); --            mac_mii_connection.mii_rx_d
		m_rx_en       : in  std_logic                     := '0';             --                              .mii_rx_dv
		m_rx_err      : in  std_logic                     := '0';             --                              .mii_rx_err
		m_tx_d        : out std_logic_vector(3 downto 0);                     --                              .mii_tx_d
		m_tx_en       : out std_logic;                                        --                              .mii_tx_en
		m_tx_err      : out std_logic;                                        --                              .mii_tx_err
		ff_rx_clk     : in  std_logic                     := '0';             --      receive_clock_connection.clk
		ff_tx_clk     : in  std_logic                     := '0';             --     transmit_clock_connection.clk
		ff_rx_data    : out std_logic_vector(31 downto 0);                    --                       receive.data
		ff_rx_eop     : out std_logic;                                        --                              .endofpacket
		rx_err        : out std_logic_vector(5 downto 0);                     --                              .error
		ff_rx_mod     : out std_logic_vector(1 downto 0);                     --                              .empty
		ff_rx_rdy     : in  std_logic                     := '0';             --                              .ready
		ff_rx_sop     : out std_logic;                                        --                              .startofpacket
		ff_rx_dval    : out std_logic;                                        --                              .valid
		ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => '0'); --                      transmit.data
		ff_tx_eop     : in  std_logic                     := '0';             --                              .endofpacket
		ff_tx_err     : in  std_logic                     := '0';             --                              .error
		ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => '0'); --                              .empty
		ff_tx_rdy     : out std_logic;                                        --                              .ready
		ff_tx_sop     : in  std_logic                     := '0';             --                              .startofpacket
		ff_tx_wren    : in  std_logic                     := '0';             --                              .valid
		ff_tx_crc_fwd : in  std_logic                     := '0';             --           mac_misc_connection.ff_tx_crc_fwd
		ff_tx_septy   : out std_logic;                                        --                              .ff_tx_septy
		tx_ff_uflow   : out std_logic;                                        --                              .tx_ff_uflow
		ff_tx_a_full  : out std_logic;                                        --                              .ff_tx_a_full
		ff_tx_a_empty : out std_logic;                                        --                              .ff_tx_a_empty
		rx_err_stat   : out std_logic_vector(17 downto 0);                    --                              .rx_err_stat
		rx_frm_type   : out std_logic_vector(3 downto 0);                     --                              .rx_frm_type
		ff_rx_dsav    : out std_logic;                                        --                              .ff_rx_dsav
		ff_rx_a_full  : out std_logic;                                        --                              .ff_rx_a_full
		ff_rx_a_empty : out std_logic                                         --                              .ff_rx_a_empty
	);
end entity Ethernet;

architecture rtl of Ethernet is
	component Ethernet_0002 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			m_rx_d        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_rx_d
			m_rx_en       : in  std_logic                     := 'X';             -- mii_rx_dv
			m_rx_err      : in  std_logic                     := 'X';             -- mii_rx_err
			m_tx_d        : out std_logic_vector(3 downto 0);                     -- mii_tx_d
			m_tx_en       : out std_logic;                                        -- mii_tx_en
			m_tx_err      : out std_logic;                                        -- mii_tx_err
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component Ethernet_0002;

begin

	ethernet_inst : component Ethernet_0002
		port map (
			clk           => clk,           -- control_port_clock_connection.clk
			reset         => reset,         --              reset_connection.reset
			reg_addr      => reg_addr,      --                  control_port.address
			reg_data_out  => reg_data_out,  --                              .readdata
			reg_rd        => reg_rd,        --                              .read
			reg_data_in   => reg_data_in,   --                              .writedata
			reg_wr        => reg_wr,        --                              .write
			reg_busy      => reg_busy,      --                              .waitrequest
			tx_clk        => tx_clk,        --   pcs_mac_tx_clock_connection.clk
			rx_clk        => rx_clk,        --   pcs_mac_rx_clock_connection.clk
			set_10        => set_10,        --         mac_status_connection.set_10
			set_1000      => set_1000,      --                              .set_1000
			eth_mode      => eth_mode,      --                              .eth_mode
			ena_10        => ena_10,        --                              .ena_10
			m_rx_d        => m_rx_d,        --            mac_mii_connection.mii_rx_d
			m_rx_en       => m_rx_en,       --                              .mii_rx_dv
			m_rx_err      => m_rx_err,      --                              .mii_rx_err
			m_tx_d        => m_tx_d,        --                              .mii_tx_d
			m_tx_en       => m_tx_en,       --                              .mii_tx_en
			m_tx_err      => m_tx_err,      --                              .mii_tx_err
			ff_rx_clk     => ff_rx_clk,     --      receive_clock_connection.clk
			ff_tx_clk     => ff_tx_clk,     --     transmit_clock_connection.clk
			ff_rx_data    => ff_rx_data,    --                       receive.data
			ff_rx_eop     => ff_rx_eop,     --                              .endofpacket
			rx_err        => rx_err,        --                              .error
			ff_rx_mod     => ff_rx_mod,     --                              .empty
			ff_rx_rdy     => ff_rx_rdy,     --                              .ready
			ff_rx_sop     => ff_rx_sop,     --                              .startofpacket
			ff_rx_dval    => ff_rx_dval,    --                              .valid
			ff_tx_data    => ff_tx_data,    --                      transmit.data
			ff_tx_eop     => ff_tx_eop,     --                              .endofpacket
			ff_tx_err     => ff_tx_err,     --                              .error
			ff_tx_mod     => ff_tx_mod,     --                              .empty
			ff_tx_rdy     => ff_tx_rdy,     --                              .ready
			ff_tx_sop     => ff_tx_sop,     --                              .startofpacket
			ff_tx_wren    => ff_tx_wren,    --                              .valid
			ff_tx_crc_fwd => ff_tx_crc_fwd, --           mac_misc_connection.ff_tx_crc_fwd
			ff_tx_septy   => ff_tx_septy,   --                              .ff_tx_septy
			tx_ff_uflow   => tx_ff_uflow,   --                              .tx_ff_uflow
			ff_tx_a_full  => ff_tx_a_full,  --                              .ff_tx_a_full
			ff_tx_a_empty => ff_tx_a_empty, --                              .ff_tx_a_empty
			rx_err_stat   => rx_err_stat,   --                              .rx_err_stat
			rx_frm_type   => rx_frm_type,   --                              .rx_frm_type
			ff_rx_dsav    => ff_rx_dsav,    --                              .ff_rx_dsav
			ff_rx_a_full  => ff_rx_a_full,  --                              .ff_rx_a_full
			ff_rx_a_empty => ff_rx_a_empty  --                              .ff_rx_a_empty
		);

end architecture rtl; -- of Ethernet
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2022 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_eth_tse" version="18.1" >
-- Retrieval info: 	<generic name="deviceFamilyName" value="MAX 10" />
-- Retrieval info: 	<generic name="core_variation" value="SMALL_MAC_10_100" />
-- Retrieval info: 	<generic name="ifGMII" value="MII" />
-- Retrieval info: 	<generic name="use_mac_clken" value="false" />
-- Retrieval info: 	<generic name="enable_use_internal_fifo" value="true" />
-- Retrieval info: 	<generic name="enable_ecc" value="false" />
-- Retrieval info: 	<generic name="max_channels" value="1" />
-- Retrieval info: 	<generic name="use_misc_ports" value="true" />
-- Retrieval info: 	<generic name="transceiver_type" value="NONE" />
-- Retrieval info: 	<generic name="enable_hd_logic" value="false" />
-- Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
-- Retrieval info: 	<generic name="enable_sup_addr" value="false" />
-- Retrieval info: 	<generic name="stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ext_stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ena_hash" value="false" />
-- Retrieval info: 	<generic name="enable_shift16" value="true" />
-- Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="false" />
-- Retrieval info: 	<generic name="enable_mac_vlan" value="false" />
-- Retrieval info: 	<generic name="enable_magic_detect" value="false" />
-- Retrieval info: 	<generic name="useMDIO" value="false" />
-- Retrieval info: 	<generic name="mdio_clk_div" value="40" />
-- Retrieval info: 	<generic name="enable_ena" value="32" />
-- Retrieval info: 	<generic name="eg_addr" value="11" />
-- Retrieval info: 	<generic name="ing_addr" value="11" />
-- Retrieval info: 	<generic name="phy_identifier" value="0" />
-- Retrieval info: 	<generic name="enable_sgmii" value="false" />
-- Retrieval info: 	<generic name="export_pwrdn" value="false" />
-- Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="phyip_pll_base_data_rate" value="1250 Mbps" />
-- Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
-- Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
-- Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
-- Retrieval info: 	<generic name="XCVR_RCFG_JTAG_ENABLE" value="0" />
-- Retrieval info: 	<generic name="XCVR_SET_CAPABILITY_REG_ENABLE" value="0" />
-- Retrieval info: 	<generic name="XCVR_SET_USER_IDENTIFIER" value="0" />
-- Retrieval info: 	<generic name="XCVR_SET_CSR_SOFT_LOGIC_ENABLE" value="0" />
-- Retrieval info: 	<generic name="XCVR_SET_PRBS_SOFT_LOGIC_ENABLE" value="0" />
-- Retrieval info: 	<generic name="enable_timestamping" value="false" />
-- Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
-- Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
-- Retrieval info: 	<generic name="AUTO_DEVICE" value="10M02DCU324A6G" />
-- Retrieval info: 	<generic name="AUTO_DEVICE_SPEEDGRADE" value="6" />
-- Retrieval info: </instance>
-- IPFS_FILES : Ethernet.vho
-- RELATED_FILES: Ethernet.vhd, Ethernet_0002.v, altera_eth_tse_mac.v, altera_tse_clk_cntl.v, altera_tse_crc328checker.v, altera_tse_crc328generator.v, altera_tse_crc32ctl8.v, altera_tse_crc32galois8.v, altera_tse_gmii_io.v, altera_tse_lb_read_cntl.v, altera_tse_lb_wrt_cntl.v, altera_tse_hashing.v, altera_tse_host_control.v, altera_tse_host_control_small.v, altera_tse_mac_control.v, altera_tse_register_map.v, altera_tse_register_map_small.v, altera_tse_rx_counter_cntl.v, altera_tse_shared_mac_control.v, altera_tse_shared_register_map.v, altera_tse_tx_counter_cntl.v, altera_tse_lfsr_10.v, altera_tse_loopback_ff.v, altera_tse_altshifttaps.v, altera_tse_fifoless_mac_rx.v, altera_tse_mac_rx.v, altera_tse_fifoless_mac_tx.v, altera_tse_mac_tx.v, altera_tse_magic_detection.v, altera_tse_mdio.v, altera_tse_mdio_clk_gen.v, altera_tse_mdio_cntl.v, altera_tse_top_mdio.v, altera_tse_mii_rx_if.v, altera_tse_mii_tx_if.v, altera_tse_pipeline_base.v, altera_tse_pipeline_stage.sv, altera_tse_dpram_16x32.v, altera_tse_dpram_8x32.v, altera_tse_dpram_ecc_16x32.v, altera_tse_fifoless_retransmit_cntl.v, altera_tse_retransmit_cntl.v, altera_tse_rgmii_in1.v, altera_tse_rgmii_in4.v, altera_tse_nf_rgmii_module.v, altera_tse_rgmii_module.v, altera_tse_rgmii_out1.v, altera_tse_rgmii_out4.v, altera_tse_rx_ff.v, altera_tse_rx_min_ff.v, altera_tse_rx_ff_cntrl.v, altera_tse_rx_ff_cntrl_32.v, altera_tse_rx_ff_cntrl_32_shift16.v, altera_tse_rx_ff_length.v, altera_tse_rx_stat_extract.v, altera_tse_timing_adapter32.v, altera_tse_timing_adapter8.v, altera_tse_timing_adapter_fifo32.v, altera_tse_timing_adapter_fifo8.v, altera_tse_top_1geth.v, altera_tse_top_fifoless_1geth.v, altera_tse_top_w_fifo.v, altera_tse_top_w_fifo_10_100_1000.v, altera_tse_top_wo_fifo.v, altera_tse_top_wo_fifo_10_100_1000.v, altera_tse_top_gen_host.v, altera_tse_tx_ff.v, altera_tse_tx_min_ff.v, altera_tse_tx_ff_cntrl.v, altera_tse_tx_ff_cntrl_32.v, altera_tse_tx_ff_cntrl_32_shift16.v, altera_tse_tx_ff_length.v, altera_tse_tx_ff_read_cntl.v, altera_tse_tx_stat_extract.v, altera_eth_tse_std_synchronizer.v, altera_eth_tse_std_synchronizer_bundle.v, altera_eth_tse_ptp_std_synchronizer.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_ecc_dec_x10.v, altera_tse_ecc_enc_x10.v, altera_tse_ecc_enc_x10_wrapper.v, altera_tse_ecc_dec_x14.v, altera_tse_ecc_enc_x14.v, altera_tse_ecc_enc_x14_wrapper.v, altera_tse_ecc_dec_x2.v, altera_tse_ecc_enc_x2.v, altera_tse_ecc_enc_x2_wrapper.v, altera_tse_ecc_dec_x23.v, altera_tse_ecc_enc_x23.v, altera_tse_ecc_enc_x23_wrapper.v, altera_tse_ecc_dec_x36.v, altera_tse_ecc_enc_x36.v, altera_tse_ecc_enc_x36_wrapper.v, altera_tse_ecc_dec_x40.v, altera_tse_ecc_enc_x40.v, altera_tse_ecc_enc_x40_wrapper.v, altera_tse_ecc_dec_x30.v, altera_tse_ecc_enc_x30.v, altera_tse_ecc_enc_x30_wrapper.v, altera_tse_ecc_status_crosser.v, altera_std_synchronizer_nocut.v
