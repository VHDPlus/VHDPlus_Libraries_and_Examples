  
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all; 

      
ENTITY Camera_CSI_Example IS
PORT (
  CLK : IN STD_LOGIC
);
END Camera_CSI_Example;

ARCHITECTURE BEHAVIORAL OF Camera_CSI_Example IS
  
BEGIN
  
END BEHAVIORAL;