-- megafunction wizard: %ALTMULT_COMPLEX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altmult_complex 

-- ============================================================
-- File Name: Complex_Mult.vhd
-- Megafunction Name(s):
-- 			altmult_complex
--
-- Simulation Library Files(s):
-- 			altera_mf;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altmult_complex CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="MAX 10" IMPLEMENTATION_STYLE="AUTO" PIPELINE=4 REPRESENTATION_A="UNSIGNED" REPRESENTATION_B="UNSIGNED" WIDTH_A=16 WIDTH_B=16 WIDTH_RESULT=32 clock dataa_imag dataa_real datab_imag datab_real result_imag result_real
--VERSION_BEGIN 18.1 cbx_alt_ded_mult_y 2018:09:12:13:04:24:SJ cbx_altera_mult_add 2018:09:12:13:04:24:SJ cbx_altera_mult_add_rtl 2018:09:12:13:04:24:SJ cbx_altmult_add 2018:09:12:13:04:24:SJ cbx_altmult_complex 2018:09:12:13:04:24:SJ cbx_arriav 2018:09:12:13:04:23:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_compare 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_parallel_add 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altmult_add 3 lpm_add_sub 7 lpm_compare 1 reg 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Complex_Mult_altmult_complex_22p IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC := '0';
		 dataa_imag	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dataa_real	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 datab_imag	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 datab_real	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 result_imag	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result_real	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END Complex_Mult_altmult_complex_22p;

 ARCHITECTURE RTL OF Complex_Mult_altmult_complex_22p IS

	 SIGNAL  wire_product1_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_product2_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_product3_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 addnsub10c	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 addnsub11c	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 addnsub12c	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_dataa	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_adder1_dataa	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_adder1_datab	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_adder1_result	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_adder2_dataa	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_adder2_datab	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_adder2_result	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor1_dataa	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_subtractor1_datab	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_subtractor1_result	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_subtractor2_dataa	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor2_datab	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor2_result	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor3_w_lg_w_result_range50w51w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor3_w_lg_w_lg_w_result_range50w51w52w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor3_dataa	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor3_datab	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor3_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor3_w_result_range50w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor4_w_lg_w_result_range48w49w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_subtractor4_dataa	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor4_datab	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor4_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_subtractor4_w_result_range48w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_comparator1_w_lg_alb25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_comparator1_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_inputb_imag_range11w30w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_inputb_imag_range11w24w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_inputb_real_range8w26w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_inputb_real_range8w31w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_addnsub47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_inputb_real_range8w26w27w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_inputb_real_range8w31w32w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add1_res :	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  addnsub :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  ena	:	STD_LOGIC;
	 SIGNAL  gnd_value :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  inputa_imag :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  inputa_real :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  inputb_imag :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  inputb_real :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  product1_res :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  product2_res :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  product3_res :	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  sub1_res :	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  sub2_res :	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_w_inputb_imag_range11w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_inputb_real_range8w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 COMPONENT  altmult_add
	 GENERIC 
	 (
		ACCUM_DIRECTION	:	STRING := "ADD";
		ACCUM_SLOAD_ACLR	:	STRING := "ACLR0";
		ACCUM_SLOAD_PIPELINE_ACLR	:	STRING := "ACLR0";
		ACCUM_SLOAD_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		ACCUM_SLOAD_REGISTER	:	STRING := "CLOCK0";
		ACCUMULATOR	:	STRING := "NO";
		ADDER1_ROUNDING	:	STRING := "NO";
		ADDER3_ROUNDING	:	STRING := "NO";
		ADDNSUB1_ROUND_ACLR	:	STRING := "ACLR0";
		ADDNSUB1_ROUND_PIPELINE_ACLR	:	STRING := "ACLR0";
		ADDNSUB1_ROUND_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		ADDNSUB1_ROUND_REGISTER	:	STRING := "CLOCK0";
		ADDNSUB3_ROUND_ACLR	:	STRING := "ACLR0";
		ADDNSUB3_ROUND_PIPELINE_ACLR	:	STRING := "ACLR0";
		ADDNSUB3_ROUND_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		ADDNSUB3_ROUND_REGISTER	:	STRING := "CLOCK0";
		ADDNSUB_MULTIPLIER_ACLR1	:	STRING := "ACLR0";
		ADDNSUB_MULTIPLIER_ACLR3	:	STRING := "ACLR0";
		ADDNSUB_MULTIPLIER_PIPELINE_ACLR1	:	STRING := "ACLR0";
		ADDNSUB_MULTIPLIER_PIPELINE_ACLR3	:	STRING := "ACLR0";
		ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1	:	STRING := "CLOCK0";
		ADDNSUB_MULTIPLIER_PIPELINE_REGISTER3	:	STRING := "CLOCK0";
		ADDNSUB_MULTIPLIER_REGISTER1	:	STRING := "CLOCK0";
		ADDNSUB_MULTIPLIER_REGISTER3	:	STRING := "CLOCK0";
		CHAINOUT_ACLR	:	STRING := "ACLR0";
		CHAINOUT_ADDER	:	STRING := "NO";
		CHAINOUT_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_ROUND_ACLR	:	STRING := "ACLR0";
		CHAINOUT_ROUND_OUTPUT_ACLR	:	STRING := "ACLR0";
		CHAINOUT_ROUND_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_ROUND_PIPELINE_ACLR	:	STRING := "ACLR0";
		CHAINOUT_ROUND_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_ROUND_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_ROUNDING	:	STRING := "NO";
		CHAINOUT_SATURATE_ACLR	:	STRING := "ACLR0";
		CHAINOUT_SATURATE_OUTPUT_ACLR	:	STRING := "ACLR0";
		CHAINOUT_SATURATE_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_SATURATE_PIPELINE_ACLR	:	STRING := "ACLR0";
		CHAINOUT_SATURATE_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_SATURATE_REGISTER	:	STRING := "CLOCK0";
		CHAINOUT_SATURATION	:	STRING := "NO";
		COEF0_0	:	NATURAL := 0;
		COEF0_1	:	NATURAL := 0;
		COEF0_2	:	NATURAL := 0;
		COEF0_3	:	NATURAL := 0;
		COEF0_4	:	NATURAL := 0;
		COEF0_5	:	NATURAL := 0;
		COEF0_6	:	NATURAL := 0;
		COEF0_7	:	NATURAL := 0;
		COEF1_0	:	NATURAL := 0;
		COEF1_1	:	NATURAL := 0;
		COEF1_2	:	NATURAL := 0;
		COEF1_3	:	NATURAL := 0;
		COEF1_4	:	NATURAL := 0;
		COEF1_5	:	NATURAL := 0;
		COEF1_6	:	NATURAL := 0;
		COEF1_7	:	NATURAL := 0;
		COEF2_0	:	NATURAL := 0;
		COEF2_1	:	NATURAL := 0;
		COEF2_2	:	NATURAL := 0;
		COEF2_3	:	NATURAL := 0;
		COEF2_4	:	NATURAL := 0;
		COEF2_5	:	NATURAL := 0;
		COEF2_6	:	NATURAL := 0;
		COEF2_7	:	NATURAL := 0;
		COEF3_0	:	NATURAL := 0;
		COEF3_1	:	NATURAL := 0;
		COEF3_2	:	NATURAL := 0;
		COEF3_3	:	NATURAL := 0;
		COEF3_4	:	NATURAL := 0;
		COEF3_5	:	NATURAL := 0;
		COEF3_6	:	NATURAL := 0;
		COEF3_7	:	NATURAL := 0;
		COEFSEL0_ACLR	:	STRING := "ACLR0";
		COEFSEL0_REGISTER	:	STRING := "CLOCK0";
		COEFSEL1_ACLR	:	STRING := "ACLR0";
		COEFSEL1_REGISTER	:	STRING := "CLOCK0";
		COEFSEL2_ACLR	:	STRING := "ACLR0";
		COEFSEL2_REGISTER	:	STRING := "CLOCK0";
		COEFSEL3_ACLR	:	STRING := "ACLR0";
		COEFSEL3_REGISTER	:	STRING := "CLOCK0";
		DEDICATED_MULTIPLIER_CIRCUITRY	:	STRING := "AUTO";
		DSP_BLOCK_BALANCING	:	STRING := "Auto";
		EXTRA_LATENCY	:	NATURAL := 0;
		INPUT_ACLR_A0	:	STRING := "ACLR0";
		INPUT_ACLR_A1	:	STRING := "ACLR0";
		INPUT_ACLR_A2	:	STRING := "ACLR0";
		INPUT_ACLR_A3	:	STRING := "ACLR0";
		INPUT_ACLR_B0	:	STRING := "ACLR0";
		INPUT_ACLR_B1	:	STRING := "ACLR0";
		INPUT_ACLR_B2	:	STRING := "ACLR0";
		INPUT_ACLR_B3	:	STRING := "ACLR0";
		INPUT_ACLR_C0	:	STRING := "ACLR0";
		INPUT_REGISTER_A0	:	STRING := "CLOCK0";
		INPUT_REGISTER_A1	:	STRING := "CLOCK0";
		INPUT_REGISTER_A2	:	STRING := "CLOCK0";
		INPUT_REGISTER_A3	:	STRING := "CLOCK0";
		INPUT_REGISTER_B0	:	STRING := "CLOCK0";
		INPUT_REGISTER_B1	:	STRING := "CLOCK0";
		INPUT_REGISTER_B2	:	STRING := "CLOCK0";
		INPUT_REGISTER_B3	:	STRING := "CLOCK0";
		INPUT_REGISTER_C0	:	STRING := "CLOCK0";
		INPUT_SOURCE_A0	:	STRING := "DATAA";
		INPUT_SOURCE_A1	:	STRING := "DATAA";
		INPUT_SOURCE_A2	:	STRING := "DATAA";
		INPUT_SOURCE_A3	:	STRING := "DATAA";
		INPUT_SOURCE_B0	:	STRING := "DATAB";
		INPUT_SOURCE_B1	:	STRING := "DATAB";
		INPUT_SOURCE_B2	:	STRING := "DATAB";
		INPUT_SOURCE_B3	:	STRING := "DATAB";
		LOADCONST_VALUE	:	NATURAL := 64;
		MULT01_ROUND_ACLR	:	STRING := "ACLR0";
		MULT01_ROUND_REGISTER	:	STRING := "CLOCK0";
		MULT01_SATURATION_ACLR	:	STRING := "ACLR1";
		MULT01_SATURATION_REGISTER	:	STRING := "CLOCK0";
		MULT23_ROUND_ACLR	:	STRING := "ACLR0";
		MULT23_ROUND_REGISTER	:	STRING := "CLOCK0";
		MULT23_SATURATION_ACLR	:	STRING := "ACLR0";
		MULT23_SATURATION_REGISTER	:	STRING := "CLOCK0";
		MULTIPLIER01_ROUNDING	:	STRING := "NO";
		MULTIPLIER01_SATURATION	:	STRING := "NO";
		MULTIPLIER1_DIRECTION	:	STRING := "ADD";
		MULTIPLIER23_ROUNDING	:	STRING := "NO";
		MULTIPLIER23_SATURATION	:	STRING := "NO";
		MULTIPLIER3_DIRECTION	:	STRING := "ADD";
		MULTIPLIER_ACLR0	:	STRING := "ACLR0";
		MULTIPLIER_ACLR1	:	STRING := "ACLR0";
		MULTIPLIER_ACLR2	:	STRING := "ACLR0";
		MULTIPLIER_ACLR3	:	STRING := "ACLR0";
		MULTIPLIER_REGISTER0	:	STRING := "CLOCK0";
		MULTIPLIER_REGISTER1	:	STRING := "CLOCK0";
		MULTIPLIER_REGISTER2	:	STRING := "CLOCK0";
		MULTIPLIER_REGISTER3	:	STRING := "CLOCK0";
		NUMBER_OF_MULTIPLIERS	:	NATURAL;
		OUTPUT_ACLR	:	STRING := "ACLR0";
		OUTPUT_REGISTER	:	STRING := "CLOCK0";
		OUTPUT_ROUND_ACLR	:	STRING := "ACLR0";
		OUTPUT_ROUND_PIPELINE_ACLR	:	STRING := "ACLR0";
		OUTPUT_ROUND_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		OUTPUT_ROUND_REGISTER	:	STRING := "CLOCK0";
		OUTPUT_ROUND_TYPE	:	STRING := "NEAREST_INTEGER";
		OUTPUT_ROUNDING	:	STRING := "NO";
		OUTPUT_SATURATE_ACLR	:	STRING := "ACLR0";
		OUTPUT_SATURATE_PIPELINE_ACLR	:	STRING := "ACLR0";
		OUTPUT_SATURATE_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		OUTPUT_SATURATE_REGISTER	:	STRING := "CLOCK0";
		OUTPUT_SATURATE_TYPE	:	STRING := "ASYMMETRIC";
		OUTPUT_SATURATION	:	STRING := "NO";
		port_addnsub1	:	STRING := "PORT_CONNECTIVITY";
		port_addnsub3	:	STRING := "PORT_CONNECTIVITY";
		PORT_CHAINOUT_SAT_IS_OVERFLOW	:	STRING := "PORT_UNUSED";
		PORT_MULT0_IS_SATURATED	:	STRING := "UNUSED";
		PORT_MULT1_IS_SATURATED	:	STRING := "UNUSED";
		PORT_MULT2_IS_SATURATED	:	STRING := "UNUSED";
		PORT_MULT3_IS_SATURATED	:	STRING := "UNUSED";
		PORT_OUTPUT_IS_OVERFLOW	:	STRING := "PORT_UNUSED";
		port_signa	:	STRING := "PORT_CONNECTIVITY";
		port_signb	:	STRING := "PORT_CONNECTIVITY";
		PREADDER_DIRECTION_0	:	STRING := "ADD";
		PREADDER_DIRECTION_1	:	STRING := "ADD";
		PREADDER_DIRECTION_2	:	STRING := "ADD";
		PREADDER_DIRECTION_3	:	STRING := "ADD";
		PREADDER_MODE	:	STRING := "SIMPLE";
		REPRESENTATION_A	:	STRING := "UNSIGNED";
		REPRESENTATION_B	:	STRING := "UNSIGNED";
		ROTATE_ACLR	:	STRING := "ACLR0";
		ROTATE_OUTPUT_ACLR	:	STRING := "ACLR0";
		ROTATE_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		ROTATE_PIPELINE_ACLR	:	STRING := "ACLR0";
		ROTATE_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		ROTATE_REGISTER	:	STRING := "CLOCK0";
		SCANOUTA_ACLR	:	STRING := "ACLR0";
		SCANOUTA_REGISTER	:	STRING := "UNREGISTERED";
		SHIFT_MODE	:	STRING := "NO";
		SHIFT_RIGHT_ACLR	:	STRING := "ACLR0";
		SHIFT_RIGHT_OUTPUT_ACLR	:	STRING := "ACLR0";
		SHIFT_RIGHT_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		SHIFT_RIGHT_PIPELINE_ACLR	:	STRING := "ACLR0";
		SHIFT_RIGHT_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		SHIFT_RIGHT_REGISTER	:	STRING := "CLOCK0";
		SIGNED_ACLR_A	:	STRING := "ACLR0";
		SIGNED_ACLR_B	:	STRING := "ACLR0";
		SIGNED_PIPELINE_ACLR_A	:	STRING := "ACLR0";
		SIGNED_PIPELINE_ACLR_B	:	STRING := "ACLR0";
		SIGNED_PIPELINE_REGISTER_A	:	STRING := "CLOCK0";
		SIGNED_PIPELINE_REGISTER_B	:	STRING := "CLOCK0";
		SIGNED_REGISTER_A	:	STRING := "CLOCK0";
		SIGNED_REGISTER_B	:	STRING := "CLOCK0";
		SYSTOLIC_ACLR1	:	STRING := "ACLR0";
		SYSTOLIC_ACLR3	:	STRING := "ACLR0";
		SYSTOLIC_DELAY1	:	STRING := "UNREGISTERED";
		SYSTOLIC_DELAY3	:	STRING := "UNREGISTERED";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL;
		WIDTH_C	:	NATURAL := 22;
		WIDTH_CHAININ	:	NATURAL := 1;
		WIDTH_COEF	:	NATURAL := 18;
		WIDTH_MSB	:	NATURAL := 17;
		WIDTH_RESULT	:	NATURAL;
		WIDTH_SATURATE_SIGN	:	NATURAL := 1;
		ZERO_CHAINOUT_OUTPUT_ACLR	:	STRING := "ACLR0";
		ZERO_CHAINOUT_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		ZERO_LOOPBACK_ACLR	:	STRING := "ACLR0";
		ZERO_LOOPBACK_OUTPUT_ACLR	:	STRING := "ACLR0";
		ZERO_LOOPBACK_OUTPUT_REGISTER	:	STRING := "CLOCK0";
		ZERO_LOOPBACK_PIPELINE_ACLR	:	STRING := "ACLR0";
		ZERO_LOOPBACK_PIPELINE_REGISTER	:	STRING := "CLOCK0";
		ZERO_LOOPBACK_REGISTER	:	STRING := "CLOCK0";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altmult_add"
	 );
	 PORT
	 ( 
		accum_sload	:	IN STD_LOGIC := '0';
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		aclr2	:	IN STD_LOGIC := '0';
		aclr3	:	IN STD_LOGIC := '0';
		addnsub1	:	IN STD_LOGIC := '1';
		addnsub1_round	:	IN STD_LOGIC := '0';
		addnsub3	:	IN STD_LOGIC := '1';
		addnsub3_round	:	IN STD_LOGIC := '0';
		chainin	:	IN STD_LOGIC_VECTOR(WIDTH_CHAININ-1 DOWNTO 0) := (OTHERS => '0');
		chainout_round	:	IN STD_LOGIC := '0';
		chainout_sat_overflow	:	OUT STD_LOGIC;
		chainout_saturate	:	IN STD_LOGIC := '0';
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clock2	:	IN STD_LOGIC := '1';
		clock3	:	IN STD_LOGIC := '1';
		coefsel0	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		coefsel1	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		coefsel2	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		coefsel3	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		dataa	:	IN STD_LOGIC_VECTOR(WIDTH_A*NUMBER_OF_MULTIPLIERS-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(WIDTH_B*NUMBER_OF_MULTIPLIERS-1 DOWNTO 0) := (OTHERS => '0');
		datac	:	IN STD_LOGIC_VECTOR(WIDTH_C*NUMBER_OF_MULTIPLIERS-1 DOWNTO 0) := (OTHERS => '0');
		ena0	:	IN STD_LOGIC := '1';
		ena1	:	IN STD_LOGIC := '1';
		ena2	:	IN STD_LOGIC := '1';
		ena3	:	IN STD_LOGIC := '1';
		mult01_round	:	IN STD_LOGIC := '0';
		mult01_saturation	:	IN STD_LOGIC := '0';
		mult0_is_saturated	:	OUT STD_LOGIC;
		mult1_is_saturated	:	OUT STD_LOGIC;
		mult23_round	:	IN STD_LOGIC := '0';
		mult23_saturation	:	IN STD_LOGIC := '0';
		mult2_is_saturated	:	OUT STD_LOGIC;
		mult3_is_saturated	:	OUT STD_LOGIC;
		output_round	:	IN STD_LOGIC := '0';
		output_saturate	:	IN STD_LOGIC := '0';
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(WIDTH_RESULT-1 DOWNTO 0);
		rotate	:	IN STD_LOGIC := '0';
		scanina	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '0');
		scaninb	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '0');
		scanouta	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		scanoutb	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		shift_right	:	IN STD_LOGIC := '0';
		signa	:	IN STD_LOGIC := '0';
		signb	:	IN STD_LOGIC := '0';
		sourcea	:	IN STD_LOGIC_VECTOR(NUMBER_OF_MULTIPLIERS-1 DOWNTO 0) := (OTHERS => '0');
		sourceb	:	IN STD_LOGIC_VECTOR(NUMBER_OF_MULTIPLIERS-1 DOWNTO 0) := (OTHERS => '0');
		zero_chainout	:	IN STD_LOGIC := '0';
		zero_loopback	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_inputb_imag_range11w30w(i) <= wire_w_inputb_imag_range11w(i) AND wire_comparator1_w_lg_alb25w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_inputb_imag_range11w24w(i) <= wire_w_inputb_imag_range11w(i) AND wire_comparator1_alb;
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_inputb_real_range8w26w(i) <= wire_w_inputb_real_range8w(i) AND wire_comparator1_w_lg_alb25w(0);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_inputb_real_range8w31w(i) <= wire_w_inputb_real_range8w(i) AND wire_comparator1_alb;
	END GENERATE loop3;
	wire_w_lg_addnsub47w(0) <= NOT addnsub(0);
	loop4 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_inputb_real_range8w26w27w(i) <= wire_w_lg_w_inputb_real_range8w26w(i) OR wire_w_lg_w_inputb_imag_range11w24w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_inputb_real_range8w31w32w(i) <= wire_w_lg_w_inputb_real_range8w31w(i) OR wire_w_lg_w_inputb_imag_range11w30w(i);
	END GENERATE loop5;
	aclr <= '0';
	add1_res <= wire_adder1_result;
	addnsub <= addnsub12c;
	ena <= '1';
	gnd_value <= (OTHERS => '0');
	inputa_imag <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & dataa_imag(15 DOWNTO 0));
	inputa_real <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & dataa_real(15 DOWNTO 0));
	inputb_imag <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & datab_imag(15 DOWNTO 0));
	inputb_real <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & datab_real(15 DOWNTO 0));
	product1_res <= wire_product1_result;
	product2_res <= wire_product2_result;
	product3_res <= ( wire_subtractor3_w_lg_w_lg_w_result_range50w51w52w);
	result_imag <= wire_adder2_result(31 DOWNTO 0);
	result_real <= wire_add_sub1_result(31 DOWNTO 0);
	sub1_res <= wire_subtractor1_result;
	sub2_res <= wire_subtractor2_result;
	wire_w_inputb_imag_range11w <= inputb_imag(15 DOWNTO 0);
	wire_w_inputb_real_range8w <= inputb_real(15 DOWNTO 0);
	product1 :  altmult_add
	  GENERIC MAP (
		INPUT_ACLR_A0 => "ACLR0",
		INPUT_ACLR_B0 => "ACLR0",
		INPUT_REGISTER_A0 => "CLOCK0",
		INPUT_REGISTER_B0 => "CLOCK0",
		MULTIPLIER_REGISTER0 => "UNREGISTERED",
		NUMBER_OF_MULTIPLIERS => 1,
		OUTPUT_ACLR => "ACLR0",
		OUTPUT_REGISTER => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		REPRESENTATION_A => "UNSIGNED",
		REPRESENTATION_B => "UNSIGNED",
		WIDTH_A => 16,
		WIDTH_B => 16,
		WIDTH_RESULT => 32
	  )
	  PORT MAP ( 
		aclr0 => aclr,
		clock0 => clock,
		dataa => inputa_real(15 DOWNTO 0),
		datab => inputb_imag(15 DOWNTO 0),
		ena0 => ena,
		result => wire_product1_result
	  );
	product2 :  altmult_add
	  GENERIC MAP (
		INPUT_ACLR_A0 => "ACLR0",
		INPUT_ACLR_B0 => "ACLR0",
		INPUT_REGISTER_A0 => "CLOCK0",
		INPUT_REGISTER_B0 => "CLOCK0",
		MULTIPLIER_REGISTER0 => "UNREGISTERED",
		NUMBER_OF_MULTIPLIERS => 1,
		OUTPUT_ACLR => "ACLR0",
		OUTPUT_REGISTER => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		REPRESENTATION_A => "UNSIGNED",
		REPRESENTATION_B => "UNSIGNED",
		WIDTH_A => 16,
		WIDTH_B => 16,
		WIDTH_RESULT => 32
	  )
	  PORT MAP ( 
		aclr0 => aclr,
		clock0 => clock,
		dataa => inputa_imag(15 DOWNTO 0),
		datab => inputb_real(15 DOWNTO 0),
		ena0 => ena,
		result => wire_product2_result
	  );
	product3 :  altmult_add
	  GENERIC MAP (
		INPUT_REGISTER_A0 => "UNREGISTERED",
		INPUT_REGISTER_B0 => "UNREGISTERED",
		MULTIPLIER_REGISTER0 => "UNREGISTERED",
		NUMBER_OF_MULTIPLIERS => 1,
		OUTPUT_ACLR => "ACLR0",
		OUTPUT_REGISTER => "CLOCK0",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		REPRESENTATION_A => "UNSIGNED",
		REPRESENTATION_B => "UNSIGNED",
		WIDTH_A => 17,
		WIDTH_B => 17,
		WIDTH_RESULT => 34
	  )
	  PORT MAP ( 
		aclr0 => aclr,
		clock0 => clock,
		dataa => add1_res(16 DOWNTO 0),
		datab => sub1_res,
		ena0 => ena,
		result => wire_product3_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN addnsub10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (ena = '1') THEN addnsub10c(0) <= wire_comparator1_alb;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN addnsub11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (ena = '1') THEN addnsub11c <= addnsub10c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN addnsub12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (ena = '1') THEN addnsub12c <= addnsub11c;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_dataa <= ( sub2_res(32 DOWNTO 0));
	wire_add_sub1_datab <= ( product3_res(32 DOWNTO 0));
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_WIDTH => 33
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_add_sub1_dataa,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	wire_adder1_dataa <= ( gnd_value & inputa_real(15 DOWNTO 0));
	wire_adder1_datab <= ( gnd_value & inputa_imag(15 DOWNTO 0));
	adder1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 17
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_adder1_dataa,
		datab => wire_adder1_datab,
		result => wire_adder1_result
	  );
	wire_adder2_dataa <= ( gnd_value & product1_res);
	wire_adder2_datab <= ( gnd_value & product2_res);
	adder2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 33
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_adder2_dataa,
		datab => wire_adder2_datab,
		result => wire_adder2_result
	  );
	wire_subtractor1_dataa <= ( gnd_value & wire_w_lg_w_lg_w_inputb_real_range8w26w27w);
	wire_subtractor1_datab <= ( gnd_value & wire_w_lg_w_lg_w_inputb_real_range8w31w32w);
	subtractor1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 17
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_subtractor1_dataa,
		datab => wire_subtractor1_datab,
		result => wire_subtractor1_result
	  );
	wire_subtractor2_dataa <= ( gnd_value & product1_res);
	wire_subtractor2_datab <= ( gnd_value & product2_res);
	subtractor2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 33
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_subtractor2_dataa,
		datab => wire_subtractor2_datab,
		result => wire_subtractor2_result
	  );
	loop6 : FOR i IN 0 TO 32 GENERATE 
		wire_subtractor3_w_lg_w_result_range50w51w(i) <= wire_subtractor3_w_result_range50w(i) AND addnsub(0);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 32 GENERATE 
		wire_subtractor3_w_lg_w_lg_w_result_range50w51w52w(i) <= wire_subtractor3_w_lg_w_result_range50w51w(i) OR wire_subtractor4_w_lg_w_result_range48w49w(i);
	END GENERATE loop7;
	wire_subtractor3_dataa <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value);
	wire_subtractor3_datab <= ( wire_product3_result(33 DOWNTO 0));
	wire_subtractor3_w_result_range50w <= wire_subtractor3_result(32 DOWNTO 0);
	subtractor3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_subtractor3_dataa,
		datab => wire_subtractor3_datab,
		result => wire_subtractor3_result
	  );
	loop8 : FOR i IN 0 TO 32 GENERATE 
		wire_subtractor4_w_lg_w_result_range48w49w(i) <= wire_subtractor4_w_result_range48w(i) AND wire_w_lg_addnsub47w(0);
	END GENERATE loop8;
	wire_subtractor4_dataa <= ( gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value & gnd_value);
	wire_subtractor4_datab <= ( wire_product3_result(33 DOWNTO 0));
	wire_subtractor4_w_result_range48w <= wire_subtractor4_result(32 DOWNTO 0);
	subtractor4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => ena,
		clock => clock,
		dataa => wire_subtractor4_dataa,
		datab => wire_subtractor4_datab,
		result => wire_subtractor4_result
	  );
	wire_comparator1_w_lg_alb25w(0) <= NOT wire_comparator1_alb;
	comparator1 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		alb => wire_comparator1_alb,
		dataa => datab_real,
		datab => datab_imag
	  );

 END RTL; --Complex_Mult_altmult_complex_22p
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Complex_Mult IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa_imag		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		dataa_real		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		datab_imag		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		datab_real		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		result_imag		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		result_real		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END Complex_Mult;


ARCHITECTURE RTL OF complex_mult IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT Complex_Mult_altmult_complex_22p
	PORT (
			clock	: IN STD_LOGIC ;
			dataa_imag	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			dataa_real	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			datab_imag	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			datab_real	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			result_imag	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			result_real	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result_imag    <= sub_wire0(31 DOWNTO 0);
	result_real    <= sub_wire1(31 DOWNTO 0);

	Complex_Mult_altmult_complex_22p_component : Complex_Mult_altmult_complex_22p
	PORT MAP (
		clock => clock,
		dataa_imag => dataa_imag,
		dataa_real => dataa_real,
		datab_imag => datab_imag,
		datab_real => datab_real,
		result_imag => sub_wire0,
		result_real => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: IMPLEMENTATION_STYLE STRING "AUTO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX 10"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "4"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "UNSIGNED"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "UNSIGNED"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa_imag 0 0 16 0 INPUT NODEFVAL "dataa_imag[15..0]"
-- Retrieval info: USED_PORT: dataa_real 0 0 16 0 INPUT NODEFVAL "dataa_real[15..0]"
-- Retrieval info: USED_PORT: datab_imag 0 0 16 0 INPUT NODEFVAL "datab_imag[15..0]"
-- Retrieval info: USED_PORT: datab_real 0 0 16 0 INPUT NODEFVAL "datab_real[15..0]"
-- Retrieval info: USED_PORT: result_imag 0 0 32 0 OUTPUT NODEFVAL "result_imag[31..0]"
-- Retrieval info: USED_PORT: result_real 0 0 32 0 OUTPUT NODEFVAL "result_real[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa_imag 0 0 16 0 dataa_imag 0 0 16 0
-- Retrieval info: CONNECT: @dataa_real 0 0 16 0 dataa_real 0 0 16 0
-- Retrieval info: CONNECT: @datab_imag 0 0 16 0 datab_imag 0 0 16 0
-- Retrieval info: CONNECT: @datab_real 0 0 16 0 datab_real 0 0 16 0
-- Retrieval info: CONNECT: result_imag 0 0 32 0 @result_imag 0 0 32 0
-- Retrieval info: CONNECT: result_real 0 0 32 0 @result_real 0 0 32 0
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: lpm
