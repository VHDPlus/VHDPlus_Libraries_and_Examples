
module LogicAnalyzer (
	acq_clk,
	acq_data_in,
	acq_trigger_in);	

	input		acq_clk;
	input	[31:0]	acq_data_in;
	input	[0:0]	acq_trigger_in;
endmodule
